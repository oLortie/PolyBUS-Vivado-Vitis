----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06/26/2021 04:45:52 PM
-- Design Name: 
-- Module Name: PolyBUS_package - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

package PolyBUS_package is
    
    ----------------------------------------------
    -- Respiration 0.25 Hz
    ----------------------------------------------
    type table_forme_respi is array (integer range 0 to 399) of std_logic_vector(11 downto 0);
    constant mem_respi025Hz : table_forme_respi := (
    -- 
    x"7FF",
    x"820",
    x"840",
    x"860",
    x"880",
    x"8A0",
    x"8C0",
    x"8E0",
    x"900",
    x"920",
    x"940",
    x"960",
    x"97F",
    x"99F",
    x"9BE",
    x"9DE",
    x"9FD",
    x"A1C",
    x"A3B",
    x"A5A",
    x"A78",
    x"A97",
    x"AB5",
    x"AD3",
    x"AF1",
    x"B0F",
    x"B2D",
    x"B4A",
    x"B67",
    x"B84",
    x"BA1",
    x"BBE",
    x"BDA",
    x"BF6",
    x"C12",
    x"C2D",
    x"C49",
    x"C64",
    x"C7F",
    x"C99",
    x"CB3",
    x"CCD",
    x"CE7",
    x"D00",
    x"D19",
    x"D31",
    x"D4A",
    x"D62",
    x"D79",
    x"D91",
    x"DA8",
    x"DBE",
    x"DD4",
    x"DEA",
    x"E00",
    x"E15",
    x"E29",
    x"E3E",
    x"E52",
    x"E65",
    x"E78",
    x"E8B",
    x"E9D",
    x"EAF",
    x"EC1",
    x"ED2",
    x"EE2",
    x"EF2",
    x"F02",
    x"F11",
    x"F20",
    x"F2F",
    x"F3C",
    x"F4A",
    x"F57",
    x"F63",
    x"F70",
    x"F7B",
    x"F86",
    x"F91",
    x"F9B",
    x"FA5",
    x"FAE",
    x"FB7",
    x"FBF",
    x"FC7",
    x"FCE",
    x"FD5",
    x"FDB",
    x"FE1",
    x"FE6",
    x"FEB",
    x"FEF",
    x"FF3",
    x"FF6",
    x"FF9",
    x"FFB",
    x"FFD",
    x"FFE",
    x"FFF",
    x"FFF",
    x"FFF",
    x"FFE",
    x"FFD",
    x"FFB",
    x"FF9",
    x"FF6",
    x"FF3",
    x"FEF",
    x"FEB",
    x"FE6",
    x"FE1",
    x"FDB",
    x"FD5",
    x"FCE",
    x"FC7",
    x"FBF",
    x"FB7",
    x"FAE",
    x"FA5",
    x"F9B",
    x"F91",
    x"F86",
    x"F7B",
    x"F70",
    x"F63",
    x"F57",
    x"F4A",
    x"F3C",
    x"F2F",
    x"F20",
    x"F11",
    x"F02",
    x"EF2",
    x"EE2",
    x"ED2",
    x"EC1",
    x"EAF",
    x"E9D",
    x"E8B",
    x"E78",
    x"E65",
    x"E52",
    x"E3E",
    x"E29",
    x"E15",
    x"E00",
    x"DEA",
    x"DD4",
    x"DBE",
    x"DA8",
    x"D91",
    x"D79",
    x"D62",
    x"D4A",
    x"D31",
    x"D19",
    x"D00",
    x"CE7",
    x"CCD",
    x"CB3",
    x"C99",
    x"C7F",
    x"C64",
    x"C49",
    x"C2D",
    x"C12",
    x"BF6",
    x"BDA",
    x"BBE",
    x"BA1",
    x"B84",
    x"B67",
    x"B4A",
    x"B2D",
    x"B0F",
    x"AF1",
    x"AD3",
    x"AB5",
    x"A97",
    x"A78",
    x"A5A",
    x"A3B",
    x"A1C",
    x"9FD",
    x"9DE",
    x"9BE",
    x"99F",
    x"97F",
    x"960",
    x"940",
    x"920",
    x"900",
    x"8E0",
    x"8C0",
    x"8A0",
    x"880",
    x"860",
    x"840",
    x"820",
    x"7FF",
    x"7DF",
    x"7BF",
    x"79F",
    x"77F",
    x"75F",
    x"73F",
    x"71F",
    x"6FF",
    x"6DF",
    x"6BF",
    x"69F",
    x"680",
    x"660",
    x"641",
    x"621",
    x"602",
    x"5E3",
    x"5C4",
    x"5A5",
    x"587",
    x"568",
    x"54A",
    x"52C",
    x"50E",
    x"4F0",
    x"4D2",
    x"4B5",
    x"497",
    x"47A",
    x"45E",
    x"441",
    x"425",
    x"409",
    x"3ED",
    x"3D1",
    x"3B6",
    x"39B",
    x"380",
    x"366",
    x"34C",
    x"332",
    x"318",
    x"2FF",
    x"2E6",
    x"2CD",
    x"2B5",
    x"29D",
    x"286",
    x"26E",
    x"257",
    x"241",
    x"22B",
    x"215",
    x"1FF",
    x"1EA",
    x"1D5",
    x"1C1",
    x"1AD",
    x"19A",
    x"187",
    x"174",
    x"162",
    x"150",
    x"13E",
    x"12D",
    x"11D",
    x"10D",
    x"0FD",
    x"0EE",
    x"0DF",
    x"0D0",
    x"0C2",
    x"0B5",
    x"0A8",
    x"09B",
    x"08F",
    x"084",
    x"079",
    x"06E",
    x"064",
    x"05A",
    x"051",
    x"048",
    x"040",
    x"038",
    x"031",
    x"02A",
    x"024",
    x"01E",
    x"019",
    x"014",
    x"010",
    x"00C",
    x"009",
    x"006",
    x"004",
    x"002",
    x"001",
    x"000",
    x"000",
    x"000",
    x"001",
    x"002",
    x"004",
    x"006",
    x"009",
    x"00C",
    x"010",
    x"014",
    x"019",
    x"01E",
    x"024",
    x"02A",
    x"031",
    x"038",
    x"040",
    x"048",
    x"051",
    x"05A",
    x"064",
    x"06E",
    x"079",
    x"084",
    x"08F",
    x"09B",
    x"0A8",
    x"0B5",
    x"0C2",
    x"0D0",
    x"0DF",
    x"0EE",
    x"0FD",
    x"10D",
    x"11D",
    x"12D",
    x"13E",
    x"150",
    x"162",
    x"174",
    x"187",
    x"19A",
    x"1AD",
    x"1C1",
    x"1D5",
    x"1EA",
    x"1FF",
    x"215",
    x"22B",
    x"241",
    x"257",
    x"26E",
    x"286",
    x"29D",
    x"2B5",
    x"2CD",
    x"2E6",
    x"2FF",
    x"318",
    x"332",
    x"34C",
    x"366",
    x"380",
    x"39B",
    x"3B6",
    x"3D1",
    x"3ED",
    x"409",
    x"425",
    x"441",
    x"45E",
    x"47A",
    x"497",
    x"4B5",
    x"4D2",
    x"4F0",
    x"50E",
    x"52C",
    x"54A",
    x"568",
    x"587",
    x"5A5",
    x"5C4",
    x"5E3",
    x"602",
    x"621",
    x"641",
    x"660",
    x"680",
    x"69F",
    x"6BF",
    x"6DF",
    x"6FF",
    x"71F",
    x"73F",
    x"75F",
    x"77F",
    x"79F",
    x"7BF",
    x"7DF" 
    -- 
    );
    
    -----------------------------------------------
    -- Respiration 0.5 Hz
    -----------------------------------------------
    type table_forme_respi2 is array (integer range 0 to 199) of std_logic_vector(11 downto 0);
    constant mem_respi05Hz : table_forme_respi2 := (
    x"7FF",
    x"840",
    x"880",
    x"8C0",
    x"900",
    x"940",
    x"97F",
    x"9BE",
    x"9FD",
    x"A3B",
    x"A78",
    x"AB5",
    x"AF1",
    x"B2D",
    x"B67",
    x"BA1",
    x"BDA",
    x"C12",
    x"C49",
    x"C7F",
    x"CB3",
    x"CE7",
    x"D19",
    x"D4A",
    x"D79",
    x"DA8",
    x"DD4",
    x"E00",
    x"E29",
    x"E52",
    x"E78",
    x"E9D",
    x"EC1",
    x"EE2",
    x"F02",
    x"F20",
    x"F3C",
    x"F57",
    x"F70",
    x"F86",
    x"F9B",
    x"FAE",
    x"FBF",
    x"FCE",
    x"FDB",
    x"FE6",
    x"FEF",
    x"FF6",
    x"FFB",
    x"FFE",
    x"FFF",
    x"FFE",
    x"FFB",
    x"FF6",
    x"FEF",
    x"FE6",
    x"FDB",
    x"FCE",
    x"FBF",
    x"FAE",
    x"F9B",
    x"F86",
    x"F70",
    x"F57",
    x"F3C",
    x"F20",
    x"F02",
    x"EE2",
    x"EC1",
    x"E9D",
    x"E78",
    x"E52",
    x"E29",
    x"E00",
    x"DD4",
    x"DA8",
    x"D79",
    x"D4A",
    x"D19",
    x"CE7",
    x"CB3",
    x"C7F",
    x"C49",
    x"C12",
    x"BDA",
    x"BA1",
    x"B67",
    x"B2D",
    x"AF1",
    x"AB5",
    x"A78",
    x"A3B",
    x"9FD",
    x"9BE",
    x"97F",
    x"940",
    x"900",
    x"8C0",
    x"880",
    x"840",
    x"7FF",
    x"7BF",
    x"77F",
    x"73F",
    x"6FF",
    x"6BF",
    x"680",
    x"641",
    x"602",
    x"5C4",
    x"587",
    x"54A",
    x"50E",
    x"4D2",
    x"497",
    x"45E",
    x"425",
    x"3ED",
    x"3B6",
    x"380",
    x"34C",
    x"318",
    x"2E6",
    x"2B5",
    x"286",
    x"257",
    x"22B",
    x"1FF",
    x"1D5",
    x"1AD",
    x"187",
    x"162",
    x"13E",
    x"11D",
    x"0FD",
    x"0DF",
    x"0C2",
    x"0A8",
    x"08F",
    x"079",
    x"064",
    x"051",
    x"040",
    x"031",
    x"024",
    x"019",
    x"010",
    x"009",
    x"004",
    x"001",
    x"000",
    x"001",
    x"004",
    x"009",
    x"010",
    x"019",
    x"024",
    x"031",
    x"040",
    x"051",
    x"064",
    x"079",
    x"08F",
    x"0A8",
    x"0C2",
    x"0DF",
    x"0FD",
    x"11D",
    x"13E",
    x"162",
    x"187",
    x"1AD",
    x"1D5",
    x"1FF",
    x"22B",
    x"257",
    x"286",
    x"2B5",
    x"2E6",
    x"318",
    x"34C",
    x"380",
    x"3B6",
    x"3ED",
    x"425",
    x"45E",
    x"497",
    x"4D2",
    x"50E",
    x"54A",
    x"587",
    x"5C4",
    x"602",
    x"641",
    x"680",
    x"6BF",
    x"6FF",
    x"73F",
    x"77F",
    x"7BF"
    );
    
    ----------------------------------------------
    -- Pression sanguine 120/80
    ----------------------------------------------
    type table_forme_pre is array (integer range 0 to 99) of std_logic_vector(11 downto 0);
    constant mem_pre12080 : table_forme_pre := (
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"001",
    x"002",
    x"005",
    x"00C",
    x"018",
    x"02E",
    x"055",
    x"095",
    x"0F9",
    x"18D",
    x"25E",
    x"372",
    x"4CB",
    x"65E",
    x"814",
    x"9CC",
    x"B5A",
    x"C94",
    x"D54",
    x"D86",
    x"D28",
    x"C4E",
    x"B1B",
    x"9BE",
    x"865",
    x"739",
    x"654",
    x"5C6",
    x"590",
    x"5A8",
    x"5FD",
    x"67E",
    x"715",
    x"7B0",
    x"83F",
    x"8B3",
    x"904",
    x"92A",
    x"921",
    x"8EA",
    x"887",
    x"7FE",
    x"757",
    x"69B",
    x"5D3",
    x"508",
    x"442",
    x"388",
    x"2DF",
    x"249",
    x"1C8",
    x"15D",
    x"105",
    x"0BF",
    x"089",
    x"061",
    x"043",
    x"02D",
    x"01E",
    x"013",
    x"00C",
    x"007",
    x"004",
    x"002",
    x"001",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000"
    );
    
    --------------------------------------------
    -- Pression 130/80
    --------------------------------------------
    constant mem_pre13080 : table_forme_pre := (
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"001",
    x"002",
    x"006",
    x"00D",
    x"01A",
    x"032",
    x"05C",
    x"0A1",
    x"10E",
    x"1AF",
    x"290",
    x"3BC",
    x"531",
    x"6E5",
    x"8C0",
    x"A9B",
    x"C4A",
    x"D9D",
    x"E6C",
    x"EA0",
    x"E38",
    x"D48",
    x"BF7",
    x"A76",
    x"8F8",
    x"7A9",
    x"6A7",
    x"600",
    x"5B6",
    x"5C0",
    x"60C",
    x"686",
    x"71A",
    x"7B2",
    x"840",
    x"8B4",
    x"904",
    x"92A",
    x"921",
    x"8EA",
    x"887",
    x"7FE",
    x"757",
    x"69B",
    x"5D3",
    x"508",
    x"442",
    x"388",
    x"2DF",
    x"249",
    x"1C8",
    x"15D",
    x"105",
    x"0BF",
    x"089",
    x"061",
    x"043",
    x"02D",
    x"01E",
    x"013",
    x"00C",
    x"007",
    x"004",
    x"002",
    x"001",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"001"
    );

    
    ----------------------------------------------
    -- Pouls 70BPM
    ----------------------------------------------
    type table_forme_pouls is array (integer range 0 to 85) of std_logic_vector(11 downto 0);
    constant mem_pouls70 : table_forme_pouls := (
    x"187",
    x"1CF",
    x"29D",
    x"3DD",
    x"57C",
    x"762",
    x"96E",
    x"B7B",
    x"D66",
    x"EFA",
    x"FF0",
    x"FFF",
    x"EE8",
    x"CBD",
    x"9BD",
    x"627",
    x"245",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"097",
    x"26F",
    x"372",
    x"39B",
    x"31F",
    x"230",
    x"103",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"013",
    x"081",
    x"0C4",
    x"0CE",
    x"0A9",
    x"06A",
    x"028",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"004",
    x"01F",
    x"034",
    x"040",
    x"046",
    x"048",
    x"04A",
    x"04C",
    x"04F",
    x"053",
    x"059",
    x"05F",
    x"065",
    x"06A",
    x"06D",
    x"06D",
    x"06B",
    x"067",
    x"061",
    x"05A",
    x"051",
    x"046",
    x"03A",
    x"02D",
    x"01E",
    x"00D",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000"
    );
    
    ---------------------------------------------
    -- Pouls 85 BPM
    ---------------------------------------------
    type table_forme_pouls2 is array (integer range 0 to 70) of std_logic_vector(11 downto 0);
    constant mem_pouls85 : table_forme_pouls2 := (
    x"093",
    x"0EF",
    x"1F3",
    x"383",
    x"582",
    x"7CB",
    x"A2D",
    x"C78",
    x"E71",
    x"FBD",
    x"FFF",
    x"EE5",
    x"C8A",
    x"93F",
    x"557",
    x"140",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"184",
    x"31C",
    x"3B3",
    x"372",
    x"299",
    x"16A",
    x"027",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"068",
    x"0AE",
    x"0B7",
    x"086",
    x"037",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"017",
    x"025",
    x"02F",
    x"036",
    x"03B",
    x"03D",
    x"03D",
    x"03A",
    x"033",
    x"029",
    x"01A",
    x"00A",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000",
    x"000"
    );
    
    ----------------------------------------------
    -- Perspiration 1
    ----------------------------------------------
    type table_forme_persp is array (integer range 0 to 99) of std_logic_vector(11 downto 0);
    constant mem_persp1 : table_forme_persp := (
    x"8A3",
    x"8B2",
    x"8C0",
    x"8CC",
    x"8CC",
    x"8C2",
    x"8B7",
    x"8AC",
    x"8A2",
    x"897",
    x"85B",
    x"81F",
    x"7E3",
    x"7A7",
    x"76B",
    x"757",
    x"743",
    x"733",
    x"733",
    x"733",
    x"767",
    x"79C",
    x"7D1",
    x"805",
    x"83A",
    x"80C",
    x"7DE",
    x"7B1",
    x"783",
    x"755",
    x"78B",
    x"7C1",
    x"7F7",
    x"82D",
    x"862",
    x"82F",
    x"7FC",
    x"7C8",
    x"795",
    x"762",
    x"743",
    x"733",
    x"733",
    x"733",
    x"733",
    x"75D",
    x"787",
    x"7B2",
    x"7DC",
    x"806",
    x"7E9",
    x"7CB",
    x"7AE",
    x"791",
    x"774",
    x"775",
    x"776",
    x"777",
    x"779",
    x"77A",
    x"797",
    x"7B4",
    x"7D1",
    x"7EF",
    x"80C",
    x"83B",
    x"86A",
    x"899",
    x"8C8",
    x"8CC",
    x"8CC",
    x"8CC",
    x"8CC",
    x"8CC",
    x"8CC",
    x"8B8",
    x"8A3",
    x"88E",
    x"879",
    x"865",
    x"836",
    x"807",
    x"7D9",
    x"7AA",
    x"77B",
    x"79F",
    x"7C3",
    x"7E7",
    x"80A",
    x"82E",
    x"846",
    x"85D",
    x"874",
    x"88C",
    x"8A3",
    x"8CC",
    x"8CC",
    x"8CC",
    x"8CC",
    x"8CC"
    );
    
    --------------------------------------------
    -- Perspiration 2
    --------------------------------------------
    constant mem_persp2 : table_forme_persp := (
    x"B10",
    x"B18",
    x"B1F",
    x"B26",
    x"B2D",
    x"B5D",
    x"B8D",
    x"BBC",
    x"BEC",
    x"C1C",
    x"BF7",
    x"BD2",
    x"BAD",
    x"B88",
    x"B63",
    x"B29",
    x"AEF",
    x"AB5",
    x"A7B",
    x"A41",
    x"A15",
    x"A14",
    x"A14",
    x"A14",
    x"A14",
    x"A33",
    x"A52",
    x"A71",
    x"A8F",
    x"AAE",
    x"A92",
    x"A75",
    x"A58",
    x"A3B",
    x"A1E",
    x"A5C",
    x"A99",
    x"AD7",
    x"B14",
    x"B52",
    x"B90",
    x"BCD",
    x"C0B",
    x"C49",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C43",
    x"C35",
    x"C27",
    x"C19",
    x"C0B",
    x"C2B",
    x"C4B",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C51",
    x"C27",
    x"BFE",
    x"BD4",
    x"BAA",
    x"B80",
    x"B8C",
    x"B97",
    x"BA3",
    x"BAF",
    x"BBA",
    x"BB2",
    x"BAA",
    x"BA1",
    x"B99",
    x"B91",
    x"B65",
    x"B39",
    x"B0D",
    x"AE1",
    x"AB6",
    x"AD9",
    x"AFC",
    x"B20",
    x"B43",
    x"B66"
    );
    
end package;
